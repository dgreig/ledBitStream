----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:40:57 07/08/2014 
-- Design Name: 
-- Module Name:    headerFile - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity headerFile is
end headerFile;

architecture Behavioral of headerFile is
constant dataBitSize: integer := 4079; -- # of bits received from pc (512bytes/510)
--constant allOnes: std_logic_vector (dataBitSize downto 0) := x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
--whiteconstant allOnes: std_logic_vector (dataBitSize downto 0) := x"5555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555";
--constant allOnes: std_logic_vector (dataBitSize downto 0) := x"000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055000055";
constant allOnes: std_logic_vector (dataBitSize downto 0) := x"202020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020002020202020202020202020202020202020202020202020202020202020202020202020202020202020002020202020202020202020202020";
--constant allOnes: std_logic_vector (dataBitSize downto 0) := x"5500000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000020000000202000";
--constant allOnes: std_logic_vector (dataBitSize downto 0) := x"202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020202020";
--constant allOnes: std_logic_vector (dataBitSize downto 0) := x"1010101000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000000000101010101010101000000000";
begin


end Behavioral;

